module one_c(a,b,c);
input a;
input b;
output reg  c;
always @ ( a or b or c)
 
endmodule
