module two_b_b(enable,d, y);
input enable;
input d;
output y;
assign y = d;
assign y = !d;
endmodule
