module one_a ( a,b,c);
input a;
input b;
output c;
assign c = a&b;
endmodule

